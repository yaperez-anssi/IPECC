--
--  Copyright (C) 2023 - This file is part of IPECC project
--
--  Authors:
--      Karim KHALFALLAH <karim.khalfallah@ssi.gouv.fr>
--      Ryad BENADJILA <ryadbenadjila@gmail.com>
--
--  Contributors:
--      Adrian THILLARD
--      Emmanuel PROUFF
--
--  This software is licensed under GPL v2 license.
--  See LICENSE file at the root folder of the project.
--

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package ecc_customize is
	-- **********************************
	-- Start of: user-editable parameters
	-- **********************************
	-- Please refer to the in-file documentation of parameters below (after the
	-- package specification), where parameters are described in the same order
	-- as they appear hereafter.
	constant nn : positive := 528;
	constant nn_dynamic : boolean := TRUE;
	type techno_type is (spartan6, virtex6, series7, ultrascale, ialtera, asic);
	constant techno : techno_type := series7; -- set a 'techno_type' value
	-- ------------------------------
	-- Performance related parameters
	-- ------------------------------
	-- multwidth is only used if 'techno' = 'asic'
	-- (otherwise its value has no meaning and can be ignored)
	constant multwidth : positive := 32; -- 32 seems fair for an ASIC default
	constant nbmult : positive range 1 to 2 := 2;
	-- parameter nbdsp below is range-constrained because it must be >=2
	constant nbdsp : positive range 2 to positive'high := 6;
	constant sramlat : positive range 1 to 2 := 1;
	constant async : boolean := TRUE;
	-- -------------------------------------------------------------
	-- Side-channel countermeasures & HW security related parameters
	-- -------------------------------------------------------------
	constant hwsecure : boolean := TRUE; -- TRUE = highly secure, FALSE = highly not
	-- hwsecure replaces the old 'debug' mode (hwsecure = TRUE <=> debug = FALSE)
	constant blinding : integer := 96; -- 96 seems fair for size of blinding rnd
	constant shuffle : boolean := TRUE; -- memory shuffling
	type shuftype is (none, linear, permute_lgnb, permute_limbs);
	constant shuffle_type : shuftype := permute_lgnb; -- set a 'shuftype' value
	constant zremask : integer := 4; -- quite arbitrary but quite often too
	-- -----------------------
	-- TRNG related parameters
	-- -----------------------
	constant notrng : boolean := TRUE; -- set to TRUE for simu, to FALSE for syn
	constant nbtrng : positive := 4;
	constant trngta : natural range 1 to 4095 := 32;
	constant trng_ramsz_raw : positive := 4; -- in kB
	constant trng_ramsz_axi : positive := 4; -- in kB
	constant trng_ramsz_efp : positive := 4; -- in kB
	constant trng_ramsz_crv : positive := 4; -- in kB
	constant trng_ramsz_shf : positive := 16; -- in kB
	-- -------------
	-- Miscellaneous
	-- -------------
	constant axi32or64 : natural := 32; -- 32 or 64 only allowed values
	constant nblargenb : positive := 32;  -- Change these two parameters only if
	constant nbopcodes : positive := 512; -- |you really know what you're doing.
	-- --------------------------
	-- Simulation-only parameters
	-- --------------------------
	constant simvecfile : string := "/tmp/ecc_vec_in.txt";
	constant simkb : natural range 0 to natural'high := 0; -- if 0 then ignored
	constant simlogfile : string := "/tmp/ecc.log";
	constant simxyshuflogfile : string := "/tmp/ecc_xyshuf.log";
	constant simtrngfile : string := "/tmp/random.txt";
	-- ********************************
	-- End of: user-editable parameters
	-- ********************************
end package ecc_customize;




--                         ******************************
--                         *      DOCUMENTATION OF      *
--                         *      ABOVE PARAMETERS      *
--                         ******************************

-- ============================================================================
-- NAME
--       'nn'
--
-- DEFINITION
--       Main security parameter.
--
-- TYPE/VALUE
--       Integer. No limit except that of the hardware ressources available
--       in your target/die-area.
--
-- DESCRIPTION
--       Defines the size in bit of large numbers implied in cryptographic
--       computations: the prime number p of course which defines the field
--       on which the elliptic curve is based on, the curve parameters a, b,
--       q of the curve, the point coordinates XP & YP of the base point, and
--       all intermediate variables used during computations.
--       Note: the order q of the curve can be greater than p (by a quantity
--       that, according to Hasse theorem, may be up to twice the square root
--       of p) therefore the value of 'nn' should be chosen as max(size of p,
--       size of q). Refer for instance to [Hankerson, Menezes, Vanstone,
--       "Elliptic Curve Cryptography", Springer 2004, p. 82, theorem 3.7],
--       or the Wikipedia article "Hasse's theorem on elliptic curves"
--       https://en.wikipedia.org/wiki/Hasse%27s_theorem_on_elliptic_curves.
--
-- SEE ALSO
--       'nn_dynamic'
--
-- ============================================================================
-- NAME
--       'nn_dynamic'
--
-- DEFINITION
--       Option to set the "dynamic prime size" feature.
--
-- TYPE/VALUE
--       Boolean (true or false).
--
-- DESCRIPTION
--       When this option is set to TRUE, it becomes possible for software
--       driver to dynamically set the security parameter, meaning the value
--       of 'nn' can be modified at runtime. This is done by writing register
--       W_PRIME_SIZE. The value statically set to 'nn' in the present file
--       then becomes the maximum value allowed at runtime. Hardware enforces
--       verification of this and, in case the condition that the value set
--       by software is greater than 'nn', raises an error flag in main status
--       register (R_STATUS) and freezes operations until a correct value
--       is set again by software.
--
--       When the option it set to FALSE, software cannot modify value of 'nn'
--       at runtime, and only cares the value set of 'nn' in the present file.
--       The advantage of setting this option to FALSE when the feature is
--       not considered useful for your own design is to save logic.
--
--       The advantage of setting this option to TRUE, when you need for your
--       own application to be able modify the security parameter at runtime,
--       is to increase performances (latency and throughput) whenever a
--       smaller value of 'nn' can be chosen.
--
-- SEE ALSO
--       'nn'
--
-- ============================================================================
-- NAME
--       'techno'
--
-- DEFINITION
--       Defines the technology (ASIC vs FPGA) you wish to target and, in the
--       FPGA case, the vendor/part.
--
-- TYPE/VALUE
--       Enumerate. Choices are between:
--         - 'series7', 'spartan6', 'ultrascale' for ARM/Xilinx FPGAs
--         - 'ialtera' for Intel-Altera FPGAs
--         - 'asic' if you're designing an ASIC or a system-on-a-chip
--
-- DESCRIPTION
--       This parameter mainly impacts the instanciation of the pipelined chain
--       of multipliers-accumulators (aka "MACC" in ASICs and "DSP blocks" in
--       FPGAs) inside each Montgomery multiplier, as this is almost the only
--       hardware feature that needs to be "black-box" instanciated in the
--       design (as opposed to inferred by synthesizer from behavorial VHDL).
--
-- SEE ALSO
--       'multwidth'
--
-- ============================================================================
-- NAME
--       'multwidth'
--
-- DEFINITION
--       Only used if 'techno' = asic, and in this case designates the size
--       of limbs in which large numbers are split and are accessible into/
--       from the memory of large numbers.
--
-- TYPE/VALUE
--       Integer. No limit a priori but you should obviously consider the
--       possible loss of performance of a multiplier which inputs would
--       become too large in your specific technological node.
--       Default of 32 seemed fair for a multiplier hardwired in an ASIC.
--
-- DESCRIPTION
--       This is the size (bitwidth) of the input operands to the multipliers
--       in the design. For sake of architectural simplicity, it is hence also
--       the bitwidth of the limbs in which large cryptographic numbers are
--       split, buffered & processed in arithmetic operations inside the IP.
--       If your design targets an FPGA, 'multwidth' is ignored and the size of
--       the limbs is given by parameter 'ww' instead (not customizable and
--       automatically set by the RTL).
--       - In an ASIC, there is obviously no predefined size for the multiplier
--         you wish to use in your design, unless your founder/standard-cell
--         library imposes you one. Therefore the designer can tweak this
--         parameter to set the area and performance of multipliers that
--         will be inferred in the hardware.
--       - In FPGA circuits, the multiplier-accumulators, which are called
--         "DSP blocks", already exist ("hard-coded") and cannot accept any
--         size of operands on their inputs. For instance the 7-series family
--         of FPGA from ARM-Xilinx offers the DSP48E1 primitive which is a
--         25x18 signed multiplier driving a(n also signed) result on 48 bits.
--         The 5 bit difference (48 - (25 + 18)) means that 5 extra bits are
--         present in the accumulator part of the DSP block to allow 32 output
--         terms of the DSP block to be added together (or added to the output
--         of neighbouring DSP blocks) without an overflow incurring. The
--         DSP blocks are performing to their best when they are instanciated
--         as a chain (aka in a pipeline) because there exist dedicated fast
--         physical connexions on both inputs and outputs of neighbouring pairs
--         of DSP blocks that bypass the general-purpose routing fabric of the
--         circuit, thus possibly incurring very high pipeline frequencies.
--         This is the architectural choice made within the IP for implementing
--         multiplications of large numbers that are required to carry on
--         Montgomery multiplications (c.f source file mm_ndsp.vhd).
--         Similarly, in the Spartan-6 family, also from ARM-Xilinx, the
--         DSP48A1 primitive allows signed 18x18 multiplications and an accumu-
--         lated output of 48 bits.
--         In Intel-Altera FPGAs such as Arrias & Stratix the DSP blocks can
--         be configured in 3 different ways: 9x9, 18x18 and 27x27, with an
--         accumulation on up to 64 bits.
--
--       The size of the limbs of large numbers manipulated in the IP (hence
--       also the size of the inputs to the multipliers) is denoted 'ww' (for
--       word's width) and is set statically (meaning at compilation/synthesis
--       time) by function 'set_ww' of package ecc_utils (file ecc_utils.vhd):
--
--         - if you have set 'techno' = asic, value of 'ww' is set to the same
--           value as 'multwidth'
--         - if target technology is an FPGA one, 'ww' is set according to the
--           'techno' parameter:
--             - for ARM-Xilinx FPGAs, 'ww' is set to 16.
--               Note: the reason for this number is that Xilinx DSP blocks
--               being either SIGNED 25x18 multipliers (in 7-series & ultra-
--               scale) or SIGNED 18x18 multipliers (in Spartan-6) multipliers,
--               only 17 bits are actually available when doing unsigned
--               arithmetics (which is what we need when splitting large
--               multiplications into smaller ones performed on limbs).
--               The MSBit is necessarily tied to a logic 0.
--               For sake of number readability when simulating the IP, the
--               value of 16 was chosen instead of 17, which should not incur
--               a significant difference in the final area nor the performance
--               of the design.
--               However if you really want to scrimp and save to the maximum,
--               you can tweak 'set_ww' function to return 17 instead of 16.
--             - for Intel-Altera FPGAs, 'ww' is set to 27. This is a peremptory
--               choice that you can also modify to a default 9 or 18 by editing
--               the code.
--
--       Note: in any of the cases described above, the VHDL code in mm_ndsp.vhd
--       performs a simple static test in order to enforce that the number of
--       chained/pipelined multiplier-accumulators cannot create an overflow on
--       the output result of the chain. The dynamic on the ouput value of the
--       chain is simply given by (2 x ww + ln2(ndsp)) where ndsp is the number
--       of multiplier-accumulator blocks in the chain (and 'ww' as defined pre-
--       viously) so the test merely consists in ensuring that this quantity
--       does not exceed the max accumulation available in accumulators of the
--       target technology.
--       (For instance in 7-series parts, DSP blocks have a 48 bit accumulator,
--       hence the maximum number of such blocks when tiled in a pipeline chain
--       is given by (2 x 16) + ln2(ndsp) = 48, which yields a huge number
--       (65536) that cannot be reached physically on one single die.
--       On the other hand, if you're targeting an ASIC and your multipliers
--       are 32x32 with an accumulator of let say 68 bit, you may only thread
--       16 MACC per Montgomery multiplier, which will usually do the job but
--       won't fit the needs of an application targeting a 521 bit security
--       (521 bit is the maximum security you may find in standardized crypto
--       protocols based on elliptic curves in 2023).
--       The numerical examples we've seen just above show you that in most
--       cases you won't have to worry about 'ww' and 'multwidth' parameters.
--
-- SEE ALSO
--       'nbdsp'
--
-- ============================================================================
-- NAME
--       'nbmult'
--
-- DEFINITION
--       Number of Montgomery multipliers instanciated in the IP.
--
-- TYPE/VALUE
--       Integer which should be kept small (default being 2)
--
-- DESCRIPTION
--       The number of Montgomery multipliers in the IP should be dictated by
--       the maximum Montgomery multiplications (aka REDC operation) that
--       can be simultaneously carried out when performing point operations
--       on a curve, that is considering one possible set of formulae for
--       point addition, point subtraction, and point doubling, among all
--       the different ones which are available from state-of-the-art.
--       In IPECC we use the so-called CoZ formulae which are available
--       in the jacobian projective representation of points. This set
--       of formulae is made possible when the points that need be added
--       do share the same Z coordinate. CoZ formulae were introduced
--       in [N. Meloni, "New point addition formulae for ECC applications",
--       2007]. A comprehensive survey can be found in [M. Rivain, "Fast and
--       Regular Algorithms for Scalar Multiplication over Elliptic Curves",
--       2011].
--       From the purely algorithmic/software point of view, CoZ formulae
--       reduce rouhgly by half the number of REDC operations needed to
--       complete one point addition, as compared to formulae that were
--       existing so far (e.g [Cohen, Miyaji, Ono, "Efficient elliptic curve
--       exponentiation using mixed coordinates", 1998]). Obviously in
--       hardware this is a matter of area/speed trade-off, however the
--       gain can be estimated by stating that the same computation speed
--       can be obtained as compared to a non-CoZ implementation with only
--       half the number of Montgomery multipliers instanciated in the hardware.
--       In IPECC by default only 2 REDC operators are instanciated in the
--       design (this is block mm_ndsp, c.f source file mm_ndsp.vhd). This is
--       the maximum number of Montgomery multiplications that it is possible
--       to carry out in parallel due to the dependency that exists between
--       intermediate variables in the CoZ formulae.
--       This means that setting 'nbmult' to a value more than 2 for your design
--       would simply increase - quite significantly - its surface, without
--       improving the speed of curve computations at all. Normally you don't
--       want to do that. On the other hand, if for any particular reason
--       you're considering choosing another set of formulae for your specific
--       design, then you may also consider tweaking parameter 'nbmult'.
--       Note that the set of formulae is implemented in software in IPECC
--       (using a custom assembly language) and can be easily edited/
--       modified. Visit the page "Explicit-Formulas Database" of website
--       hyperelliptic.org for a comprehensive description of elliptic curve
--       formulae, with a comparison of their performances.
--
-- ============================================================================
-- NAME
--       'nbdsp'
--
-- DEFINITION
--       Number of MACC/DSP blocks per Montgomery multipliers
--
-- TYPE/VALUE
--       Integer greater or equal to 2
--
-- DESCRIPTION
--       This parameter directly influences the performance of the IP by
--       allowing you to control the area/speed trade-off in the Montgomery
--       multipliers.
--       Obviously the more there are MACC/DSP blocks in each Montgomery
--       multiplier, the less it will take for them to carry out a complete
--       REDC operation.
--       Note however that the "speed vs nbdsp" relation is linear only
--       in a specific range of the 'nbdsp' parameter, a range which can
--       sometimes turn to be quite small - meaning that past a specific
--       threeshold (that is dependent mainly on the values of 'nn' and 'ww')
--       the computation speed obviously will plateau however hard you try
--       and increase parameter 'nbdsp' (actually it may even decrease due to
--       the fact that the excess of MACC/DSP blocks will increase the time
--       for data to go through the chain without increasing the number of
--       usefull multiplications per clock cycle).
--       The table below gives the duration in microseconds of one REDC
--       operation for 'nn' = 256 in 'techno' = 'asic', for different values
--       of the parameter 'ww' (which in the case of asic matches 'multwidth')
--       and different values of the 'nbdsp' parameter.
--       The mm_ndsp block is assumed to run at 300 MHz.
--
--            \ nbdsp |   2    3    4    5    6     8     10   12   13
--          ww \      |
--        ------------+--------------------------------------------------
--           8        | 12.8  9    7.8  6.7  6.1   5.5    5    4.5  4.5
--          16        |  4.3  3.3  3    2.7  2.4   2.4    2.2  2.2
--          32        |  1.8  1.4  1.4
--          64        |   .9   .8   .9
--
--       Note that the static value of parameter 'nn' determines the maximum
--       value allowed for 'nbdsp', which matches the number of 'ww'-bit limbs
--       large numbers are made of. Function set_ndsp in package ecc_pkg.vhd
--       enforces that this limit is not exceeded, it is used to compute the
--       value of a parameter called 'ndsp' (based on 'nbdsp') which is the
--       constant actually used in the RTL code: if value of 'nbdsp' set by
--       user in present file is below the limit, then 'ndsp' = 'nbdsp', and
--       if it is greater, then ndsp is set to the limit.
--       For instance in the example above and with 'ww' = 16, the limit to
--       'nbdsp' is 17, therefore any value for 'nbdsp' above 17 will be
--       ignored and replaced by 17. Now the table above also tells us that
--       17 is already a suboptimal value for 'nbdsp', and that you'd probably
--       better set 'nbdsp' = 10 instead.
--
-- ============================================================================
-- NAME
--       'sramlat'
--
-- DEFINITION
--       Read latency for all the blocks of SRAM memory used in the IP
--
-- TYPE/VALUE
--       Integer, with only values 1 or 2 allowed.
--
-- DESCRIPTION
--       All SRAM blocks instanciated in the IP are purely synchronous and
--       have the same latency when accessed in read mode, which can be either
--       1 or 2 clock cycles, as defined by this parameter.
--       Choosing 2 instead of 1 simply means trying to increase the maximum
--       frequency at the cost of an extra layer of flip-flops on the output
--       data bus. This can be of interest in particular in FPGAs as the
--       SRAM blocks are natively provided with this extra layer of registers
--       inside the block itself, which is why synthesizer will most probably
--       infer to use these internal registers instead of consuming flip-flops
--       from the general logic fabric. Hence for an FPGA technology you pro-
--       bably want to set this parameter to 2.
--
-- ============================================================================
-- NAME
--       'async'
--
-- DEFINITION
--       If TRUE, the Montgomery multipliers in the design will reside in
--       a specific clock-domain (independent of the rest of the IP).
--
-- TYPE/VALUE
--       Boolean (true or false).
--
-- DESCRIPTION
--       This is an attempt at a "globally asynchronous / locally synchronous"
--       feature in the IP.
--       The Montgomery multiplication is notoriously the most costful operation
--       in asymetric cryptography algorithms, so the purpose of this option is
--       to allow the designer to isolate the Montgomery multipliers in their
--       own specific clock-domain that can thus be optimized as regards to
--       timing considerations.
--       You may try to:
--         - increase the frequency of that specific clock domain without
--           stressing the backend tools on the remaining parts of the circuit,
--           as they are less impacting on performances
--         - perform timing optimization solely on this clock domain as it
--           is the one that deserves the highest optimization effort.
--       Obviously the two aspects are related and should be analyzed together.
--
--       Depending on the value of 'async' paramter, the clock-domains in the IP
--       are as follows:
--         - if 'async' = FALSE, then there is only one clock-domain and the IP
--           is totally synchronous to the same clock, which thus also happens
--           to be the clock of the AXI-interconnect the IP is connected to.
--         - if 'async' = TRUE, then there are two clock-domains in the IP.
--           One clock-domain is the one in which data transfers are made on
--           the AXI-interconnect and all arithmetic operationsa except REDC
--           are also carried out.
--           The second clock-domain is the one of the REDC operators (Montgo-
--           mery multipliers).
--           In this case the usual synchronization issues at the crossing
--           of the domains are resolved in two differents ways:
--             - for control signals a layer of two or three resynchroniozation
--               flip-flops is used
--             - for data signals, we use the fact that most FPGA families offer
--               asynchronous dual-port memories to push data in one clock
--               domain and pull them in another without having to worry about
--               synchronization issues (possible metastability in the read
--               clock-domain that would be due to asynchronicity with write
--               clock will be gone by the time data are actually read).
--           If you're targeting an ASIC, you should first check the availabi-
--           lity of single dual port (asynchronous) memories in your technolo-
--           gical library.
--
--       Note having solely one clock-domain may be penalizing in FPGAs if the
--       SoC and interconnect (the IP is connected to) imposes you to run at a
--       low frequency. Values such as 100 or 150 MHz are typically found in
--       SoC-FPGA ecosystems however this is not the highest frequency by far
--       that you can hope the Montgomery multipliers to run at. Actually 200
--       MHz should be seen as the minimum target on the 28-nm node FPGAs such
--       as the ARM-Xilinx 7-series family or Ithe ntel-Altera Stratix V family.
--
--       If 'async' is set to FALSE, then the unique input clock to the IP is
--       the 's_axi_aclk' input port on top-level 'ecc' entity.
--       If 'async' is set to TRUE, 's_axi_aclk' is still the primary clock
--       input, and the dedicated clock to the REDC operators must be driven
--       on 'clkmm' input port of the IP top-level.
--
-- ============================================================================
-- NAME
--       'hwsecure'
--
-- DEFINITION
--       To choose between 'HW secure mode' versus 'HW unsecure mode' of the IP.
--
--       In a nutshell, Hw unsecure mode means any tampering with the IP is made
--       easy to the software driver. On the contrary HW secure mode means
--       hardware security is at its max.
--
--       Setting 'hwsecure' to FALSE is very dangerous in a product and should
--       not apply to production purposes, as this mode allows software driver
--       to tamper in any possible way with the IP, making it possible for each
--       security feature and countermeasure to be disengaged at runtime at the
--       software initiative.
--
--       Setting 'hwsecure' to TRUE is what you wish if you're targeting pro-
--       duction mode and you aim at disposing of a true hardware secure
--       element for your application.
--
-- TYPE/VALUE
--       Boolean, true or false.
--
-- DESCRIPTION
--       The IP can be used in two different modes which are exclusive of one
--       another: either the IP is configured in HW secure mode or it is confi-
--       gured in HW unsecure/Side-Channel analysis mode (HW unsecure mode for
--       short). This configuration is static and can’t be modified at runtime.
--       Setting 'hwsecure' to FALSE naturally means setting the IP in the
--       HW unsecure mode, and in HW secure mode otherwise.
--
--       HW unsecure mode means that interacting with the IP through software
--       driver is made very permissive, so as to allow pre-production analysis
--       of the IP and of its side-channel leakages. Software driver can then
--       tamper freely with almost any security feature implemented in the IP.
--
--       In HW unsecure mode, software-driver can:
--         - read or write the value of any large number in memory, at any time
--         - insert breakpoints into microcode to interrupt scalar multiplica-
--           tion and perform step by step execution (e.g to allow time iso-
--           lation of a specific part of [k]P computation for clean, reduced-
--           noise side-channel measurement)
--         - specify a precise time in the course of [k]P computation where to
--           activate or deactivate the trigger signal driven out of the IP
--           (this is 'dbgtrigger' output port of top-level entity 'ecc').
--           Use cases for the external out trigger feature include oscilloscope
--           input-trigger activation and EM injection probe setting-off.
--           This feature is clock-cycle accurate
--         - bypass the TRNG and force use of deterministic numbers instead of
--           random ones
--         - access internal memory array of the TRNG raw random bit FIFO, in
--           order to perform entropy quality assessment
--         - modify the content of the microcode memory to implement and
--           evaluate different curve formulae or different countermeasures.
--         - enable or disable almost any of the countermeasures.
--
--       In HW secure mode:
--         - the only large numbers software driver is allowed to WRITE in
--           memory are the first eight ones (large number address 0 to 7).
--           These are: prime number p, curve parameters a, b and q, scalar k
--           and base point coordinates XP & YP
--         - the only large numbers software driver is allowed to READ from
--           memory are:
--             - the two coordinates of the result point (these are
--               x_{[k]P} and y_{[k]P} in affine representation) which are avai-
--               lable for read at the same address as XP and YP are respecti-
--               vely available for write)
--             - the one-shot random masking token that the IP uses to whiten
--               the [k]P result coordinates. Software driver is required to
--               read that number before ordering any [k]P computation, other-
--               wise it won't be able to obtain the plain (unmasked) value of
--               the [k]P result coordinates.
--         - breakpoints do not exist (control logic & data paths are pruned
--           at synthesis time)
--         - outside trigger does not exit (control logic & data paths are
--           pruned at synthesis time).
--         - TRNG cannot be bypassed, nor random values be forced, nor random
--           values be read by software (control logic and read data paths are
--           pruned at synthesis time)
--         - microcode memory cannot be modified (content is fixed at syn-
--           thesis time and write data path to memory is pruned).
--         - Interactions between software driver and IP are strongly res-
--           tricted. Whenever software issues a command that requires
--           computation from the IP, it can no longer issues any command
--           before that computation is totally carried out and completed.
--         - The choice made by the hardware designer at synthesis time on
--           the following 3 options : 'blinding', 'shuffle', and 'zremask'
--           can only be modified by the software driver if it increases
--           the level of security. For instance, if 'blinding' is 0 in
--           ecc_customize.vhd, it means software driver will still be able
--           to program [k]P computations with blinding. On the other hand,
--           if 'blinding' > 0, then software driver won't be able to suppress
--           blinding at runtime. Same applies to 'shuffle', and same applies
--           to 'zremask' (the 'shuffle' parameter however behaves a bit dif-
--           ferently in the sense that if 'shuffle' = FALSE statically in
--           ecc_customize.vhd, then it can't be activated at runtime, see
--           below description of parameter 'shuffle').
--           The idea behind the three parameters named 'blinding', 'zremask'
--           and 'shuffle' (along with 'shuffle_type') is to allow the hardware
--           designer, to lock the corresponding countermeasure as always
--           applicable to each [k]P computation, and it is important to keep
--           in mind that these locks are effective only if you also set at
--           the same time parameter 'hwsecure' to TRUE.
--           Setting 'hwsecure' parameter to FALSE instead would actually
--           maintain the possibility to engage each of these countermeasures,
--           but at the discretion of the software driver and on a [k]P-compu-
--           tation per [k]P-computation basis.
--           Note that 'blinding', 'shuffle' & 'zremask' features are not the
--           only side-channel countermeasures provided with the IP, but only
--           those that you can choose to statically hardlock. This is because
--           they are the most performance costly.
--
--       To sum-up:
--
--         - If you intend to use the IP in a security application such as a
--       Secure Element, a Hardware Security Module or if you entend to
--       integrate it as hardware accelerator inside a general purpose SoC,
--       choose FALSE.
--
--         - If you intend to use the IP for an academic/research purpose,
--       to evaluate the side-channel resistance of the IP on a specific
--       target, or during the preproduction phase of your product, choose
--       TRUE (in the latter case, you may consider to "logic-lock" all
--       the portion of the design that will remain when you eventually
--       turn the parameter to FALSE and send it to foundry).
--
-- REMARK
-- 
--       'hwsecure' has replaced paremeter 'debug' starting from v1.4.6,
--       with the equivalence hwsecure = not debug (hwsecure = TRUE is
--       equivalent to old 'debug' parameter = FALSE, and hwsecure = FALSE
--       is equivalent to old 'debug' parameter = TRUE).
--
--       Some parts of the code have kept the debug_/_debug/_debug_/_dbg/
--       or _DBG token in a few signal names, driver API functions, etc,
--       but it doesn't change anything to their definition. When you see
--       "debug" in the code/comments, it means "HW unsecure".
--
-- SEE ALSO
--       'blinding', 'shuffle', 'zremask'
--
-- ============================================================================
-- NAME
--       'blinding'
--
-- DEFINITION
--       This parameter is used to statically activate (and configure), or
--       statically deactivate the blinding side-channel countermeasure.
--
-- TYPE/VALUE
--       Integer.
--       0 means disable, otherwise any strictly positive number will set
--       the bit size of the blinding number.
--       Default is 96.
--
-- DESCRIPTION
--       When non null, 'blinding' gives the bit size of the random number
--       "alpha" used to randomize the original scalar "k" set by software,
--        according to equation:
--
--                             k' = k + (alpha x q)
--
--       where "q" designates the order of the elliptic curve.
--
--       The rule of thumb is to set a bitwidth of approx. 96 for 'nn' = 256.
--       Hardware enforces that the size be smaller than 'nn' (either the
--       static value when 'nn_dynamic' = FALSE, or the runtime dynamic one
--       when 'nn_dynamic' = TRUE).
--
--       Setting 0 instead will keep the blinding countermeasure available but
--       solely as an option that software can decide to set or not to set at
--       each [k]P computation.
--
-- IMPORTANT NOTE:
--       Setting a non-0 value to 'blinding' only makes sense if you also set
--       'hwsecure' to TRUE.
--       If you set 'hwsecure' to FALSE, the value set for 'blinding' won't make
--       a difference as software driver will then be considered legitimate
--       in modifying the blinding settings at runtime, including the possi-
--       bility to completely disable blinding.
--
-- SEE ALSO
--       'hwsecure', 'shuffle', 'zremask'
--
-- ============================================================================
-- NAME
--       'shuffle'
--
-- DEFINITION
--       This parameter is used to statically activate or statically deactivate
--       the shuffling side-channel countermeasure.
--
-- TYPE/VALUE
--       Boolean (true or false)
--       Default is true.
--
-- DESCRIPTION
--       The purpose of the shuffling countermeasure is to break the relation
--       between large numbers and the address in the physical memory they are
--       read from during sensitive computations.
--
--       When set to TRUE, 'shuffle' parameter activates the random shuffling of
--       the complete memory storing large cryptographic numbers between the
--       processing of each bit of the scalar. This countermeasure thwarts the
--       attacks aimed at guessing which intermediate variables are manipulated
--       inside point addition formulae by use of their address's physical
--       leakage. As memory shuffling removes the relation between addresses
--       and values of the aforementioned variables, these attacks become
--       infeasible - or at least much difficult to be carried out.
--
--       Set to TRUE if you want the shuffling of large numbers' memory to be
--       activated at each [k]P computation (memory is shuffled inbetween the
--       processing of two consecutive bits of the scalar). The method used to
--       to shuffle the memory is then defined as per parameter 'shuffle_type'.
--
--       Setting FALSE instead to 'shuffle' parameter will keep the counter-
--       measure available (if parameter 'shuffle_type' is different than
--       'none', see below) but solely as an option that software can decide
--       to use or not to use at each [k]P computation.
--
--       In any case, the choice of the shuffling method is static as only one
--       can be implemented at synthesis time, among 'linear', 'permute_lgnb'
--       and 'permute_limbs' (see parameter 'shuffle_type' below).
--
--       Setting 'shuffle' to TRUE only makes sense if you also set 'hwsecure'
--       to TRUE. If you set 'hwsecure' to FALSE, the value set for 'shuffle'
--       won't make a difference, as software driver will then be considered
--       legitimate in modifying the shuffle settings at runtime, including
--       the possibility to completely disable it.
--
-- SEE ALSO
--       'shuffle_type', 'hwsecure', 'blinding', 'zremask'
--
-- ============================================================================
-- NAME
--       'shuffle_type'
--
-- DEFINITION
--       Defines the way large numbers' memory is shuffled.
--       This parameter is relevant even if 'shuffle' = FALSE, because
--       it defines what will be synthesized (and hence instanciated) in
--       the hardware.
--       For instance setting:
--          - 'shuffle' = FALSE
--       together with:
--          - 'shuffle_type' = linear
--       means that a linear shuffling method will be synthesized, however
--       shuffling won't be forced; instead it will be applied only if
--       software driver enables shuffling (with register W_SHUFFLE).
--
-- TYPE/VALUE
--       One of 'linear', 'permute_lgnb', 'permute_limbs' or 'none'.
--       Default is 'permute_lgnb'.
--
-- DESCRIPTION
--
--       The three available methods of shuffling correspond to a compromise
--       between implementation complexity & perf. cost on one side, and
--       efficiency as a side-channel countermeasure on the other.
--
--       The 'linear' method is simple to implement and should incur almost
--       no performance penalty at all (neither in surface nor on speed).
--       The 'permute_limbs' method should quite damage the speed performance,
--       and is probably "overkill". Besides, as discussed below, as it requires
--       an SRAM block memory to store the address indirection, it is possible
--       that its gain might not be real in terms of side-channel resistance.
--       It is also expected to consume large quantities of randomness.
--       The 'permute_lgnb' method offers an intermediate solution, both in
--       terms of surface and speed, which makes it probably the best solution
--       (which is why it was set as the default choice).
--
--       The description below first covers the two "extreme" methods ('linear'
--       and 'permute_limbs'), 'permute_lgnb' being explained last.
--
--       'linear':
--
--          Shuffling will consist in drawing a random mask and applying it
--          linearly (xor) to the read address of each data word to determine
--          the target (shuffled) write address. Therefore when the counter-
--          measure is activated the memory is physically duplicated inside
--          the IP and a flip/flop mechanism is used to ensure consistency
--          of the transfer of one version of the memory into its newly shuf-
--          fled version.
--          The address here designates the address of *limbs* inside the
--          large numbers' memory. Hence limbs of the large numbers are what
--          is shuffled here, meaning that each one of the 'nblargenb' large
--          numbers stored in memory will have its 'ww'-bit limbs scattered
--          all accross the memory array, however their addresses will keep
--          a linear relation between them.
--          The number of possible permutations in this case is not very
--          important. For instace for 'nn' = 256 and 'ww' = 16 (and assuming
--          the default value of 32 for 'nblargenb', the address of a 'ww'-bit
--          limb in memory will be of 10 bits, which makes it a total of 2**10
--          (1024) different possible permutations (this should be compared to
--          the 1024! ways of permutating a memory array of 1024-words, which
--          is what is offered by the 'permute_limbs' method).
--
--       'permute_limbs':
--
--          This method consists in permutating the large numbers' memory using
--          the Fisher-Yates algorithm.
--          Generally speaking, the Fisher-Yates algorithm is used to randomly
--          generate any permutation of an n-element set 'a' among the total n!
--          possibilities of doing so. The algorithm is very simple and consists
--          in scanning the n items (for instance in the range 'i' from 'n - 1'
--          downto 0), generating for each step 'i' a random number j in [0..i],
--          and swapping the items of the set 'a' in positions 'i' & 'j' (noted
--          a[i] <-> a[j]).
--          The difference between the 'permute_limbs' & 'permute_lgnb' methods
--          of shuffling is that in the former the Fisher-Yates algorithm is ap-
--          plied on limbs, while in the latter it is applied on whole large
--          numbers.
--          Hence in the 'permute_limbs' method, many performance aspects of
--          the implementation are expected to decrease: [k]P computation time
--          mmight probably increase a lot, and an important throughout will
--          probably required for randomness. Furthermore, and this is probably
--          the worst, it is obvious that a second SRAM block memory is made
--          necessary in the implementation in order to store the definition of
--          the permutation at any time. Well, the presence of an SRAM memory
--          in order to store the large numbers was already a drawback in itself
--          (from the perspective of side-channels (*)) that the shuffling
--          countermeasure was intended at mitigating in the first place.
--          Using another SRAM block to store the permutation (i.e the address
--          translation table) might therefore not be the more judicious to
--          do so. That's the reason for the option 'permute_lgnb' described
--          hereafter. The advantage of the 'linear' option is also that it won't
--          be synthesized but in logic gates, not memory.
--          (Finally the option 'permute_limbs' was kept in the source code to
--          allow experiments).
--
--              (*) For instance in FPGAs all physical memories have the same
--                  size (typically 32 kbit) therefore the physical leakage
--                  occuring while reading a large number from its RAM block
--                  is expected to be the same as the one that would occur when
--                  reading the randomized address from another RAM block.
--                  Power consumption as well as EM emission in digital cir-
--                  cuits is proportional to the capacitive load of nets,
--                  which are quite important in memory physical layouts.
--          
--       'permute_lgnb':
--
--          Here "lgnb" stands for large numbers, meaning the Fisher-Yates algo-
--          rithm is used to permutate whole large numbers (not only their
--          limbs). Considering the default value of 32 for the number of large
--          numbers stored in memory, it is then possible to synthesize the
--          translation table as a tiny memory of 160 bits (32 words of 5 bits)
--          whose side-channel signature should be a lot weaker than the large
--          large numbers' memory, while still allowing the complete 32! permu-
--          tations (~10^35) to be equally feasible (the component named
--          'virt_to_phys_ram_async' which implements this memory describes an
--          asynchronous read memory in order to enforce this synthesis result
--          in FPGAs (in Xilinx FPGA, the translation memory could thus be
--          synthesized using only 4 LUT located in the same slice).
--
-- NOTE:
--       As opposed to 'blinding' & 'zremask', it is not possible for the
--       software driver to enable shuffling if option 'shuffle' was not
--       statically set to TRUE, nor it is possible to modify the shuffling
--       method dynamically (meaning at runtime).
--
--       If 'shuffle' = TRUE, then only one shuffling method will be synthe-
--       sized and present in the hardware, according to the value of parame-
--       ter 'shuffle_type'. If moreover 'hwsecure' = FALSE, then software
--       driver will be able to enable or disable the shuffling.
--
--       Now if 'shuffle' = FALSE, software driver won't be able to activate
--       it. This is because the hardware implementing the shuffling of memory
--       won't be present in the circuit to begin with.
-- 
-- SEE ALSO
--       'shuffle', 'nblargenb', 'hwsecure', 'blinding', 'zremask'
--
-- ============================================================================
-- NAME
--       'zremask'
--
-- DEFINITION
--       Used to enable or disable statically the periodic repetition, all
--       along the course of [k]P computation, of random re-generation of the
--       coordinates of sensitive points, using each time a new fresh random
--       value. This countermeasure is based on the so-called Jacobian projec-
--       tive representation which by definition uses 3 coordinates (X : Y : Z)
--       to characterize points on an elliptic curve, instead of two in the
--       affine (x, y) system.
--
-- TYPE/VALUE
--       Integer.
--       A value of 0 disables the countermeasure, yet software driver will
--       still be able to activate it at rutime.
--       Default value is 4 but this is quite arbitrary. You should consider
--       the performance penalty induced by the countermeasure when selecting
--       the value for this parameter (and when doing so, keep in mind that
--       the smaller the value, the bigger the performance loss) - see last
--       paragraph of section DESCRIPTION below for performance considera-
--       tions.
--
-- DESCRIPTION
--       For 'zremask' parameter, setting a non-0 integer will define a periodi-
--       city, expressed in number of bits of the scalar, at which the coordina-
--       tes of points R0 and R1 (used throughout the scalar loop to compute
--       [k]P) will be re-randomized using a fresh multiplicative random (aka
--       "Z-masking" countermeasure). Note that such a masking is always applied
--       at the beginning of the scalar loop, regardless of value set for
--       'zremask'. What you can set with 'zremask' is to force that masking to
--       happen again and periodically throughout the entire scalar loop.
--       With e.g default setting 'zremask' = 4, coordinates will be rando-
--       mized with a new fresh random every one in four bits of the scalar.
--
--       There is a 1-1 correspondence between the set of affine points
--
--                               {(x, y) : x,y \in F_p}
--
--       and the set of projective points
--
--                        {(X : Y : Z) : X,Y,Z \in F_p, Z != 0}
--
--       verifying x = X / (Z**2),  y = Y / (Z**3).
--       Hence the Z coordinate can be used as some kind of "free" variable
--       allowing us to choose between virtually an infinite number (actually
--       p - 1) of ways to represent any point on the elliptic curve. For any
--       valid representation (X : Y : Z) that belongs to the equivalence class
--       of an affine point (x, y) then for any number L in F_p \ {0}, the tri-
--       plet { (L^2).X : (L^3).Y : L.Z } belongs to the same equivalence class,
--       hence represents the same point.
--       This countermeasure has been called "Randomized projective coordina-
--       tes" in the paper that originally introduced the idea (c.f [J.-B.
--       Coron, "Resistance against Differential Power Analysis for Elliptic
--       Curve Cryptosystems", CHES'1999]). In the context of the IP we call
--       that countermeasure "Z-remasking" as the idea is to allow the user of
--       of the IP/designer of the hardware system to repeat the randomization
--       of the point representation several times inside each [k]P represen-
--       tation.
--
--       Setting 'zremask' = 0 will keep the Z-masking countermeasure available
--       but solely as an option that software can decide to set or not to set
--       at each [k]P computation.
--
--       Setting a non-0 value to 'zremask' only makes sense if you also set
--       'hwsecure' to TRUE (if you set 'hwsecure' to FALSE, the value set for
--       'zremask' won't make a difference as software driver will then be
--       considered legitimate in modifying the 'zremask' settings at runtime
--       or simply disabling it).
--
--       Note that when option 'nn_dynamic' is set to TRUE, the value set for
--       'zremask' is independent of the runtime value 'nn' can take. If for
--       instance 'zremask' = 4, re-randomization will happen every 4 bits of
--       the scalar whether 'nn' = 256 or 'nn' = 384. But while in the former
--       case it will happen 64 times throughout the whole [k]P computation,
--       it will happen 96 times in the latter.
--
--       The cost of the countermeasure is 8 REDC (8 Montgomery multiplications)
--       at each remasking, so you'd better consider the performance cost of
--       setting the countermeasure 'zremask', given that each bit of the scalar
--       already costs 16 REDC per itself in Co-Z representation (which is the
--       one used in the IP). Obviously the performance cost decreases as the
--       value of 'zremask' increases (choosing for instance 'zremask' = 1 would
--       mean randomly refreshing the point coordinates after each bit of the
--       scalar, which would dramatically increase the computation cost of the
--       [k]P operation).
--
-- SEE ALSO
--       'hwsecure'
--
-- ============================================================================
-- NAME
--       'notrng'
--
-- DEFINITION
--       Used to amputate the testbench from the TRNG HDL despcription
--       which is not fit to simulation and replace it with a file containing
--       "random" data.
--       MUST BE SET TO FALSE IN SYNTHESIS (otherwise synthesis will fail)
--       AND TO TRUE IN SIMULATION (otherwise simulation will hang).
--
-- TYPE/VALUE
--       Boolean (true or false).
--       Default is TRUE, hence fitting simulation. Change to FALSE before
--       synthesis!
--
-- DESCRIPTION
--       The HDL description of the TRNG in the IP contains a combinational
--       loop which cannot be simulated (it would hang the simulator engine
--       by creating an infinite number of simulation steps (deltas) inside
--       each physical instant). This is why you must set this parameter
--       depending on what you're doing with the IP, simulating it or synthe-
--       sizing it:
--
--         - when you're simulating, parameter 'notrng' must be set to TRUE.
--           All the ES-TRNG instances are then removed from the HDL model, as
--           well as the binary tree gathering their outputs (see below discus-
--           sion of parameter 'nbtrng'). Instead a simulation-only process is
--           instanciated that will read "random" data from the file specified
--           in parameter 'simtrngfile' (see below this parameter).
--
--         - when you're synthesizing, parameter 'notrng' must be set to FALSE.
--           The HDL model then embeds the ES-TRNG component with the combina-
--           tional loop describing the ring oscillator.
--
--       If you provided the IP with a random post-processor (again refer to
--       discussion for parameter 'nbtrng' below) it will still be part of
--       the simulation model when 'notrng' = TRUE.
--
-- WARNING
--       Vivado tool from ARM-Xilinx seems not comfortable with this parameter
--       being set to either one of "/dev/random" or "/dev/urandom" (it will
--       halt simulation from the begining).
--
-- SEE ALSO
--       'simtrngfile'
--
-- ============================================================================
-- NAME
--       'nbtrng'
--
-- DEFINITION
--       Number of TRNG primitives instanciated in parallel in the IP.
--
-- TYPE/VALUE
--       Integer which should be set according to the entropy throughput
--       required for a specific application. Default is 1.
--
-- BIBLIO
--       [Yang, Rozic, Grujic, Mentens, Verbauwhede, "ES-TRNG, A High-
--       throughput, Low-area True Random Number Generator based on Edge
--       Sampling"]
--       (https://tches.iacr.org/index.php/TCHES/article/view/7276)
--       
-- DESCRIPTION
--       The physical true random number generator used in the IP is the
--       ES-TRNG, designed at the COSIC research group of KU Leuven. It was
--       first published at the CHES'18 conference. Its architecture makes it
--       particularly suitable to FPGA designs. It has a very small footprint,
--       while still exhibiting very good throughput results.
--       Porting it to an ASIC technology should not be difficult as the
--       only FPGA-specific features that it relies on are carry propagation
--       primitives (usually used for adders and counters) which are actually
--       used in ES-TRNG as pure delay propagation lines. ASIC buffers would
--       normally fit this purpose without any problem.
--
--       We do not give here the architecture nor the design principles of
--       ES-TRNG, rather we point the reader to its online presentation paper
--       (c.f section BIBLIO above).
--
--       The way ES-TRNG is used in the IP is that exactly 'nbtrng' copies
--       of the ES-TRNG primitive are physically instanciated in the IP.
--       They operate completely independently one from the other and
--       "periodically" generate a random bit along with its strobe signal
--       (the quotation marks on word "periodically" are because each random
--       bit itself is generated after a period of accumulation of jitter
--       which is itself random, althought there is a minimum for that delay
--       which is given by parameter 'trngta' - see below).
--       The outputs of each different instances of ES-TRNG primitive are
--       gathered together using a binary routing tree that terminates with
--       a unique root output. (Althought not required, it is probably best
--       that you set a power of two for value of 'nbtrng').
--       Due to the average number of clock cycles it will take for each
--       ES-TRNG primitive to issue one random bit (this number is related to
--       'trngta' parameter, see below) congestion of the tree is not to be
--       expected unless you really set too large a value for 'nbtrng'.
--       Ideally this parameter should be set to a number such that at each
--       clock cycle, and given the frequency at which the IP main clock is
--       set, a new random bit presents itself at the root of the tree.
--       Output raw random bits are pushed into a FIFO which feeds a post-
--       processing unit.
--
--       +===============================================================+
--       | THE POST-PROCESSING UNIT IS NOT PART OF THE IPECC DESIGN AND  |
--       | SHOULD BE PROVIDED BY YOUR OWN CARE. THE ROLE OF POST-PRO-    |
--       | CESSING FUNCTION IN RANDOM APPLICATIONS IS IMPORTANT BECAUSE  |
--       | IT GUARANTEES THAT THE OUPUT OF THE RANDOM GENERATOR REMAINS  |
--       | UNPREDICTABLE TO AN ATTACKER EVEN IF SHE TAKES CONTROL OF THE |
--       | PHYSICAL ENTROPY SOURCE AND THAT THE OUTPUT OF THE PHYSICAL   |
--       | ENTROPY SOURCE BECOMES DETERMINISTIC TO HER (e.g THROUGH A    |
--       | "STUCK-AT-0" OR A "STUCK-AT-1" INVASIVE OR SEMI-INVASIVE KIND |
--       | OF ATTACK).                                                   |
--       +===============================================================+
--
--       In present release of the IP, as no postprocessing unit is provided,
--       the output port of the raw random bit FIFO is directly connected to
--       the logic that would normally extract postprocessed bits. This "logic
--       stub" allows the IP to be operational as is - that is, despite the
--       absence of postprocessing on the raw random bits - while allowing
--       to very simply plug any cryptographic logic component that you may
--       design or reuse to implement the postprocessing, provided that its
--       interfaces fit the ones we use inside the IP TRNG (which are very
--       basic).
--
--       Past the postprocessing unit, random bits are pushed one at a time
--       into one of the 4 possible target FIFOs, each serving as the entropy
--       pool for one of the 4 features/countermeasures of the IP that require
--       random data. These 4 features are:
--
--         1. the on-the-fly masking of the scalar in the AXI interface, at the
--            time it is pushed by software driver in the memory of large
--            numbers;
--         2. the NNRND instruction which IP microcode can use to generate a
--            complete random large number in the memory of large numbers;
--         3. the 4-by-4 shuffling that the IP applies to the 4 coordinates
--            XR0, YR0, XR1 and YR1 of points R0 and R1 inbetween the processing
--            of each bit of the scalar;
--         4. the shuffling countermeasure of the complete memory of large
--            numbers, when it is set and activated (see parameter 'shuffle'
--            above).
--
--       A round-robin scheduling is applied to the bits pulled from the
--       postprocessing unit to ensure that each of the 4 target FIFOs fairly
--       gets the same amount of random data as long as it is not already full.
--       Needless to say, no bit pushed in any of the 4 FIFOs gets aslo
--       pushed in any of the three others. The 4 FIFOs aare this filled
--       with completely independent random bits.
--
--       The sizes of each of the 4 target FIFOs are defined in the package
--       file ecc_trng/ecc_trng_pkg.vhd. The default sizes are functions of
--       the parameter 'nn' (directly or indirectly, as some depends on
--       parameter 'n' which in turn depends on 'nn' and 'ww'). If you need
--       to customize the amount of random data equired for each of the 4
--       features in your application, you may do it in this file.
--
--       In HW unsecure mode, diagnostic features allow you to read the
--       content of the raw random bit memory through the AXI interface in
--       order to perform statisticial tests and estimate the entropy of each
--       TRNG instances (the entropy performance of each instance directly
--       relies on its floorplan realization, therefore they won't be
--       necessarily the same for all instances).
--
--       For FPGA applications, the design rationale you should apply here
--       is that once the entropy quality s estimated good enough of one
--       instance (this is assessed using statistical tests suits such as
--       the one provided by U.S NIST or german BSI) you should "logic-lock"
--       this instance using the software feature that CAD tools provide
--       you with, preventing the instance from being re-placed or re-routed
--       elsewhere in future place-and-route runs of your circuit.
--
--       Note that the IP does not include statistical self-tests.
--
-- IMPORTANT
--       The default setting of 1 for parameter 'nbtrng' might not be sufficient
--       to your application!
--       You must perform a throughput analysis and evaluation of the randomness
--       your application specifically needs, and set, along with a properly
--       chosen 'trngta' parameter, the number of ES-TRNG instances that is fit
--       to achieve this throughput.
--       The effect of not assessing the quantity/throughput of entropy your
--       application needs is that the IP might often stall at runtime. This
--       will happen each time the IP needs to perform an operation that
--       requires a minimum amount of entropy to be properly carried out till
--       the end, and that amount is not available yet in the corresponding
--       FIFO.
--
-- SEE ALSO
--       'trngta', 'notrng'
--
-- ============================================================================
-- NAME
--       'trngta'
--
-- DEFINITION
--       Main sizing parameter of the entropy quality generated by the ES-TRNG
--       primitive.
--
-- TYPE/VALUE
--       Integer. Default is 32 but this value is quite arbitrary.
--
-- DESCRIPTION
--       The greater the value of 'trngta' is, the highest the entropy per
--       random bit is, but also the smaller the random production througput.
--       The smaller the value of 'trngta' is, the greater the throughput is,
--       but also the poorer the entropy per bit is.
--
--       The principle of ES-TRNG is the same as many other TRNG designs: a free
--       running oscillator is formed using a ring of inverters in odd number,
--       and let to run freely until a specific amount of time is passed so as
--       to consider that enough entropy has been accumulated in the phase noise
--       ("jitter" in the time domain) of the oscillator edges. Value of para-
--       meter 'trngta' exactly denotes the duration of that "free-running"
--       phase of the oscillator, expressed in number of periods of the main
--       system clock of the IP. (Remember from what was stated earlier - see
--       'async' section above -, that is clock is the one connected to the
--       input port 's_axi_aclk' of the top-level entity). The meaning of the
--       value of 'trngta' therefore depends on the frequency of that main
--       clock and it carries no sense without it.
--       When the free-running phase has passed, some very tiny logic (that can
--       fit into a very small number of FPGA LUTs) is triggered to detect the
--       first rising edge of the free oscillator. This detector samples the
--       information as to whether the sampling clock "saw" the edge of the
--       oscillator before or after its own edge, thus capturing in one bit
--       the jitter of the free-oscillator.
--
--       Only tests and measurements made on real hardware can assess that
--       number properly.
--
-- SEE ALSO
--       'nbtrng', 'notrng'
--
-- ============================================================================
-- NAME
--       'trng_ramsz_[raw|axi|efp|crv|shf]'
--
-- DEFINITION
--       These 5 parameters each set the size of one of the FIFO used to
--       buffer random numbers inside the IP before they are serviced to
--       their respective entropy clients.
--
-- TYPE/VALUE
--       All 5 parameters are integer, expressed in kilo-bytes.
--
-- DESCRIPTION
--       In terminology of AIS31 standard, parameter 'trng_ramsz_raw' is
--       related to "raw random numbers", which are random numbers directly
--       taken at the output of the physical source, before any logical
--       "post-processing". Other 4 parameters 'trng_ramsz_[axi|efp|crv|shf]
--       are related to "internal random numbers" (AIS31 terminology again),
--       which are random numbers taken at the output of the post-processing
--       operations.
--       Each of the 5 parameters is translated (this is done in package
--       ecc_trng_pkg) into an associated parameter expressing the size of
--       the same FIFO, but this time in number of elements (or "words") of
--       the corresponding FIFO's memory array. Moreover, they are ROUNDED UP
--       TO THE NEXT (OR EQUAL) POWER OF 2.
--
--         - 'trng_ramsz_raw' is translated into parameter 'raw_ram_size'.
--           Now as the raw random FIFO stores bits, we obviously have:
--
--             'raw_ram_size' = greater or equal power-of-2 of qty
--                                (  8 * 1024 * 'trng_ramsz_raw' )
--
--         - 'trng_ramsz_axi' is translated into parameter 'irn_fifo_size_axi'.
--           The FIFO of internal random nb served to ecc_axi storing ww-bit
--           words, we have:
--
--             'irn_fifo_size_axi' = greater or equal power-of-2 of qty
--                                 ( 'trng_ramsz_axi' * 1024 * 8) / ww )
--
--         - 'trng_ramsz_efp' is translated into parameter 'irn_fifo_size_efp'.
--           The FIFO of internal random nb served to ecc_fp storing ww-bit
--           words, we have:
--
--             'irn_fifo_size_efp' = greater or equal power-of-2 of qty
--                                 ( 'trng_ramsz_efp' * 1024 * 8) / ww )
-- 
--         - 'trng_ramsz_crv' is translated in parameter 'irn_fifo_size_crv'.
--           The FIFO of internal random nb served to ecc_curve storing 2-bit
--           words, we have:
--
--             'irn_fifo_size_crv' = greater or equal power-of-2 of qty
--                                 ( 'trng_ramsz_crv' * 1024 * 8) / 2 )
--
--         - 'trng_ramsz_shf' is translated into parameter 'irn_fifo_size_shf'.
--           The FIFO of internal random nb served to ecc_fp_dram_sh_* storing
--           words whose bitwidth depends on the type of shuffling algorithm
--           selected by parameter 'shuffle_type' (see that parameter and its
--           description), parameter 'irn_fifo_size_shf' is deduced from
--           'trng_ramsz_shf' through a relation similar as those above but
--           depending on the parameter 'shuffle_type' (see VHDL function
--           'set_irn_width_sh' defined in package file ecc_pkg.vhd and used
--           in ./ecc_trng/ecc_trng_pkg.vhd).
--
-- SEE ALSO
--       'nbtrng', 'notrng', 'shuffle_type'
--
-- ============================================================================
-- NAME
--       'axi32or64'
--
-- DEFINITION
--       Defines the width of the data buses of the AXI interfaces of the IP.
--       These are: the WDATA signal bus of the AXI-lite write-data channel,
--       and the RDATA signal bus of the AXI-lite read-data channel.
--
-- TYPE/VALUE
--       Integer, with only values 32 or 64 allowed.
--
-- DESCRIPTION
--       To simplify integration of the IP inside any AXI-interconnect/system-
--       on-chip (meaning: independently of whether the architecture is 32 or
--       64 bit) registers accessible by the software driver:
--
--         - are all 32-bit long (as if data buses were that of a 32-bit
--           system), WITH THE EXCEPTION OF THE TWO REGISTERS W_WRITE_DATA
--           and R_READ_DATA;
--
--         - have address aligned on 8 bytes (as if address buses were that
--           of a 64-bit system).
--
--       The size of both registers W_WRITE_DATA and R_READ_DATA depends on
--       parameter 'axi32or64':
--
--         - when the IP is configured using 'axi32or64' = 32, then W_WRITE_DATA
--           and R_READ_DATA are 32 bit long.
--           Therefore, if the AXI-interconnect the IP is connected to is 64 bit
--           then:
--
--             - when reading register R_READ_DATA, the 32 upper bits of the
--               signal bus RDATA (AXI read data channel) will be cleared
--               (zeroed) by the IP
--
--             - when writing register W_WRITE_DATA, the 32 upper bits of the
--               signal bus WDATA (AXI write data channel) will be ignored
--               by the IP.
--
--         - when the IP is configured using 'axi32or64' = 64, then W_WRITE_DATA
--           and R_READ_DATA are 64 bit long.
--           Therefore, if the AXI-interconnect the IP is connected to is
--           32 bit, then you might consider adding extra logic in between the
--           IP and the AXI-interconnect so as to:
--
--             - gather two consecutive read accesses to R_READ_DATA into one
--               64 bit read transaction to the IP and split the result into
--               two 32-bit responses to transaction initiator (CPU, memory
--               controller, bridge, etc).
--
--             - gather two consecutive write accesses to W_WRITE_DATA into
--               one 64 bit write transaction to the IP.
--
--             In both cases (read & write) software should be aware of the
--             mismatch between size of the IP AXI interface and the size of
--             the AXI interconnect, so that to enforce that transactions
--             should always be issued by pair (otherwise deadlock might occur).
--
-- IMPORTANT NOTE:
--       Experiments made on real hardware, namely Xilinx(R) Zynq(R) SoC/FPGA
--       platforms, show that is is probably better to always set parameter
--       'axi32or64' to 32. These real-hardware tests indeed showed that even
--       when the IP was connected to an AXI 64-bit interface (and despite
--       the fact that Cortex-A53 used for these tests were 64-bit cores)
--       bus transactions issued from the CPU were still 32-bit ones, thus
--       incurring data errors with an IP configured in mode 'axi32or64' = 64.
--
--       In any case, set 'axi32or64' = 64  *ONLY IF*  you are absolutely
--       sure and have characterized, in your own hardware application, the
--       property that AXI transactions emitted by the CPU when writing
--       (resp. reading) to register W_WRITE_DATA (resp. from register
--       R_READ_DATA) are 64-bit transactions and that they will never be
--       split in 32-bit transactions during their complete path through the
--       interconnect from the CPU to the IP (resp. from the IP to the CPU).
--
--       The restriction descrived above probably narrows down the utility
--       of parameter 'axi32or64', which hence might be suppressed in future
--       releases of the IP.
--
-- ============================================================================
-- NAME
--       'nblargenb'
--
-- DEFINITION
--       Number of cryptographic large numbers that inner memory of the IP
--       can buffer.
--
-- TYPE/VALUE
--       Integer. Default is 32. Obviously keep it a power of 2.
--
-- DESCRIPTION
--       Note that this is not a memory size in bytes or bits or whatever
--       absolute unity of size, this is a relative number. For instance
--       if each large number is 256 bit wide, then the size of the memory of
--       large numbers will be given by 32 x 256 bit = 8 Kbit (assuming the
--       default of 32 for parameter 'nblargenb').
--
--       The IP is basically an ALU for large numbers controlled by a hardware
--       state machine that fetches and decodes arithmetic instructions opera-
--       ting on these large numbers. An opcode format exists for such instruc-
--       tions describing in particular the address of the numbers in the
--       memory of large numbers which are to be read and/or written by each
--       instruction. Most of instructions contain 3 operands named opa, opb &
--       opc, with opa & opb being the input (read) operands & opc the output
--       (written) operand. All these fields are, in the current release of the
--       IP, 5 bit address fields pointing to a large number. This value of 5
--       bit obviously matches the size of the memory, which is made of 32
--       large numbers. The 32 default was chosen because it is the minimum
--       that we were able to fit into the set of all intermediate variables
--       involved in the computation of the scalar multiplication (the most
--       complex operation performed by the IP). To that default setting of 32
--       large numgers corresponds 5-bit fields for addresses op[abc] in the
--       instruction opcodes, which packed along other fields turned out to
--       to form a quite practical 32-bit size for the opcode words.
--
--       You can change the value of parameter 'nblargenb', but you should do
--       it with precaution. The HDL code of the IP was written all along with
--       genericity in mind, notably regards the parameters 'nblargenb' &
--       'nbopcodes' (see below) however not many simulation runs nor tests
--       were actually done with other values than the default ones (resp. 32
--       and 512). So you should change these parameters only if you really
--       know that you're doing.
--
--       Mind in particular that increasing the value of 'nblargenb' will
--       have the size of fields op[abc] in instruction opcodes obviously
--       also increase (e.g to 6 bit if you set 'nblargenb' to 64). This in
--       turn will make opcodes become larger than 32 bit.
--
-- ============================================================================
-- NAME
--       'nbopcodes'
--
-- DEFINITION
--       Size of the microcode memory of the IP, in number of instruction
--       opcodes.
--
-- TYPE/VALUE
--       Integer. Default is 512. Same as 'nblargenb' above: obviously keep it
--       a power of 2.
--
-- DESCRIPTION
--       Note that this is not a memory size in bytes or bits or whatever
--       absolute unity of size, this is a relative number. For instance
--       if size of each opcode is 32 bit wide (the default) then the
--       physical size of the microcode memory will be given by 512 x 32 bit
--       = 16 Kbit (assuming the default of 512 for parameter 'nbopcodes').
--
--       Please refer to the discussion above for parameter 'nblargenb',
--       as it also widely applies to 'nbopcodes'.
--
-- ============================================================================
-- NAME
--       'simvecfile'
--
-- DEFINITION
--       Only used in simulation.
--       Name of the input file providing input test-vector files to the
--       simulation testbench (we name this file the "input test-vector file").
--
-- TYPE/VALUE
--       Character string indicating a file path which should be accessible
--       in read mode.
--
-- DESCRIPTION
--       The format expected for the file pointed to by 'simvecfile' is the
--       exact same format as the one of the input test-vector file expected
--       by the program 'ecc-test-linux-uio' (or 'ecc-test-linux-devmem')
--       aimied at testing the real hardware (see sources in folder 'driver/').
--       Please refer to the Appendix of main documentation PDF (doc/ipecc.pdf)
--       titled "Simulating the IP".
--
--       IMPORTANT NOTE: The input test-vector file is not expected to provide
--       only entry values for the tests (curve parameters and base point coor-
--       dinates). What is meant here is that the file SHOULD ALSO contain the
--       RESULT expected for each test (e.g the coordinates of [k]P, or the
--       answer 'true' or 'false' of a boolean test). The simulation testbench
--       (or the test program of the real hardware) will submit the test input
--       data to the IP, run the expected command, then collect the result back
--       from the IP and compare it with what is provided as the expected output
--       in the input test-vector file.
--
--       Please refer to the script file <generate-tests.sage> (in folder 'sage/')
--       for a quick and easy way to generate an input test vector file. This
--       script contains a start section that includes the definition of all
--       the parameters required for the generation of tests (that you can
--       obviously customize to meet your requirements) including an online
--       textual help on each of these parameters.
--
-- ============================================================================
-- NAME
--       'simkb'
--
-- DEFINITION
--       Only used in simulation, to artificially restrict the size of a large
--       scalar.
--
-- TYPE/VALUE
--       Integer. Must be greater than or equal to 3.
--
-- DESCRIPTION
--       When 'simkb' is different from 0, then the main right-to-left loop
--       which parses the scalar bits will span only bits 0 to simkb - 1.
--       You can therefore use parameter 'simkb' as if you were truncating
--       the scalar set by software driver to its lowest 'simkb' bits, without
--       modifying your simulation testbench.
--
--       When 'simkb' is 0, then the main loop will parse all the bits of the
--       scalar.
--
-- WARNING
--       It doesn't make sense to restrict the size of the scalar (using
--       'simkb') in a simulation where blinding countermeasure is also
--       enabled, or at least simply keep in mind that the quantity of bits
--       that will be taken into account by the IP are the ones of the
--       *blinded* scalar, hence the result can bear no more logic relation
--       to the scalar as it was set initially by the software driver.
--
-- ============================================================================
-- NAME
--       'simlogfile'
--
-- DEFINITION
--       Only used in simulation. File path for the simulation trace log.
--
-- TYPE/VALUE
--       Character string indicating a file path which should be accessible
--       in write mode.
--       Default is "/tmp/ecc.log" which should be convenient (at least for
--       Unix-like systems).
--
-- DESCRIPTION
--       This is the path of the file where simulation will dump the information
--       detailing all the instructions that were executed by ecc_curve.vhd,
--       with the address of thier operands, their result, timestamp, etc.
--
--       If you provide a relative path, the place where the file will actually
--       be placed is dependent on your simulator (the default "/tmp/ecc.log"
--       was made an absolute path to avoid this). If you provide a simple file-
--       name, Vivado will likely create it in 'sim_1/behav/xsim/' in your local
--       project folder.
--
-- ============================================================================
-- NAME
--       'simtrngfile'
--
-- DEFINITION
--       Only used in simulation.
--       Name of the input file providing "random" data to the TRNG simulation
--       testbench.
--
-- TYPE/VALUE
--       Character string indicating a file path which should be accessible
--       in read mode.
--       Default is "/tmp/random.txt" is arbitrary.
--
-- DESCRIPTION
--       Format of this file is the following: each value should be an
--       unsigned decimal integer ranging from 0 to 255, with one value
--       per line.
--       Simulation will stop when it hits the end of the file.
--
--       File sim/HOWTO-random.txt gives an example of a one-liner
--       command you can use to quickly generate this file.
--
-- SEE ALSO
--       'notrng'
